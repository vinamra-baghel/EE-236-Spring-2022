Vinamra Baghel 190010070 Schottky IV Characteristics

.include schottky_BAT85.txt
.include schottky_BAT960.txt
.include Diode_1N914.txt

*Netlist
r1 in 1 100
r2 3 gnd 100
r3 1 gnd 1k
X1 1 2 BAT85
Vdr1 2 3 0

r4 in 4 100
r5 6 gnd 100
r6 4 gnd 1k
X2 4 5 BAT960
Vdr2 5 6 0

r7 in 7 100
r8 9 gnd 100
r9 7 gnd 1k
D3 7 8 1N914
Vdr3 8 9 0

Vin in gnd 0

*Analysis
.dc Vin 0 5 0.01

.control
run
set color0 = white
set color1 = black
set color2 = red
set color3 = blue
set color4 = green
set xbrushwidth = 2
plot I(Vdr1) vs V(1)-V(2) I(Vdr2) vs V(4)-V(5) I(Vdr3) vs V(7)-V(8)
*let Vd1 = V(1)-V(2)
*meas dc Vd1 find Vd1 when I(Vdr) = 1m
.endc
.end