Vinamra Baghel 190010070 CMOS Inverter Transient Characteristics

.include CMOS.txt

*Netlist
M11 out1 in dd dd cmosp L=0.4u W=60u AS=48p PS=121.6u AD=48p PD=121.6u
M12 out1 in 0 0 cmosn L=0.4u W=30u AS=24p PS=61.6u AD=24p PD=61.6u
Cl1 out1 0 0.05p

M21 out2 in dd dd cmosp L=0.4u W=60u AS=48p PS=121.6u AD=48p PD=121.6u
M22 out2 in 0 0 cmosn L=0.4u W=60u AS=48p PS=121.6u AD=48p PD=121.6u
Cl2 out2 0 0.05p

M31 out3 in dd dd cmosp L=0.4u W=30u AS=24p PS=61.6u AD=24p PD=61.6u
M32 out3 in 0 0 cmosn L=0.4u W=60u AS=48p PS=121.6u AD=48p PD=121.6u
Cl3 out3 0 0.05p

Vdd dd 0 3.3
Vin in 0 pulse(0 3.3 0 20p 20p 4n 8n 0)

*Analysis
.tran 0.01n 10n

.control
run
set color0 = white
set color1 = black
set color2 = red
set color3 = blue
set color4 = green
set color5 = orange
set xbrushwidth = 3

plot V(in) V(out1) V(out2) V(out3)

meas tran tr1 trig V(out1) val=0.1*3.3 td=0 rise=1 targ V(out1) val=0.9*3.3 td=0 rise=1
meas tran tf1 trig V(out1) val=0.9*3.3 td=0 fall=2 targ V(out1) val=0.1*3.3 td=0 fall=2

meas tran tr2 trig V(out2) val=0.1*3.3 td=0 rise=1 targ V(out2) val=0.9*3.3 td=0 rise=1
meas tran tf2 trig V(out2) val=0.9*3.3 td=0 fall=2 targ V(out2) val=0.1*3.3 td=0 fall=2

meas tran tr3 trig V(out3) val=0.1*3.3 td=0 rise=1 targ V(out3) val=0.9*3.3 td=0 rise=1
meas tran tf3 trig V(out3) val=0.9*3.3 td=0 fall=2 targ V(out3) val=0.1*3.3 td=0 fall=2

print tr1 tf1 tr2 tf2 tr3 tf3

meas tran tin when V(in)=1.65
meas tran tout1 when V(out1)=1.65
print tout1-tin
meas tran tout2 when V(out2)=1.65
print tout2-tin
meas tran tout3 when V(out3)=1.65
print tout3-tin
.endc
.end