Vinamra Baghel 190010070 IV Characteristics Part 1

.include Diode_1N914.txt
.include rn142s.txt

*Netlist
r1 in out1 100
D1 1 gnd DRN142S
Vd1 out1 1 0

r2 in out2 100
D2 2 gnd 1N914
Vd2 out2 2 0

Vin in gnd 0

*Analysis
.dc vin 0 5 0.1

.control
run
set color0 = white
set color1 = black
set color2 = red
set color3 = blue
set xbrushwidth = 3
plot I(Vd1) vs V(1) I(Vd2) vs V(2)

meas dc i11 find I(Vd1) when V(1) = 810m
meas dc i12 find I(Vd1) when V(1) = 800m
let il11 = log(abs(i11))
let il12 = log(abs(i12))
let e1 = 10m/(((273+75)/298)*26m*(il11-il12))

meas dc i21 find I(Vd2) when V(2) = 810m
meas dc i22 find I(Vd2) when V(2) = 800m
let il21 = log(abs(i21))
let il22 = log(abs(i22))
let e2 = 10m/(((273+75)/298)*26m*(il21-il22))

print e1 e2
.endc
.end