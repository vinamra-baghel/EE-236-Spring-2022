Vinamra Baghel 190010070 Schottky Bridge Rectifier

.include schottky_BAT85.txt
.include schottky_BAT960.txt

*Netlist
rl out1 out2 1k
X1 in out2 BAT85
X2 out1 in BAT85
X3 out1 gnd BAT85
X4 gnd out2 BAT85
Vin in gnd sin(0 12 50 0 0 0)

*Analysis
.tran 1u 60m

.control
run
set color0 = white
set color1 = black
set color2 = red
set color3 = blue
set xbrushwidth = 2
plot V(out2) - V(out1)
.endc
.end