Vinamra Baghel 190010070 CMOS Inverter

.include CMOS.txt

*Netlist
M11 out1 in dd dd cmosp L=0.4u W=60u AS={2*60u*0.4u} PS={2*60u+4*0.4u} AD={2*60u*0.4u} PD={2*60u+4*0.4u}
M12 out1 in 0 0 cmosn L=0.4u W=30u AS={2*30u*0.4u} PS={2*30u+4*0.4u} AD={2*30u*0.4u} PD={2*30u+4*0.4u}
Cl1 out1 0 0.05p

Vdd dd 0 3.3
Vin in 0 0

*Analysis
.dc Vin 0 3.3 0.01 Vdd 1.5 3 1.5

.control
run
set color0 = white
set color1 = black
set color2 = red
set color3 = blue
set color4 = green
set color5 = orange
set xbrushwidth = 3

let Vout1 = V(out1)[0, 330]
let Vout2 = V(out1)[331, 661]
plot Vout1 vs V(in)[0, 330] Vout2 vs V(in)[331, 661]

.endc
.end